module hello_world;

initial begin
$display("Hello World by Abhay Pawar");
#20 $finish;

end
endmodule